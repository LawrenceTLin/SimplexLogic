treat mom